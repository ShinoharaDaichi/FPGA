	component test is
		port (
			clk_clk             : in std_logic := 'X'; -- clk
			reset_reset_n       : in std_logic := 'X'; -- reset_n
			spi_0_reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component test;

	u0 : component test
		port map (
			clk_clk             => CONNECTED_TO_clk_clk,             --         clk.clk
			reset_reset_n       => CONNECTED_TO_reset_reset_n,       --       reset.reset_n
			spi_0_reset_reset_n => CONNECTED_TO_spi_0_reset_reset_n  -- spi_0_reset.reset_n
		);

