library verilog;
use verilog.vl_types.all;
entity timer_vlg_check_tst is
    port(
        hordiv          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end timer_vlg_check_tst;
