-- blinker.vhd

-- Generated using ACDS version 15.0 145

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity blinker is
	port (
		clk_clk                             : in  std_logic                    := '0';             --                          clk.clk
		led_external_connection_export      : out std_logic_vector(7 downto 0);                    --      led_external_connection.export
		switcher_external_connection_export : in  std_logic_vector(7 downto 0) := (others => '0')  -- switcher_external_connection.export
	);
end entity blinker;

architecture rtl of blinker is
	component blinker_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component blinker_led;

	component blinker_nios2_proc is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component blinker_nios2_proc;

	component blinker_onchip_memory is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(63 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(63 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(7 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component blinker_onchip_memory;

	component blinker_switcher is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component blinker_switcher;

	component blinker_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component blinker_sysid_qsys_0;

	component blinker_mm_interconnect_0 is
		port (
			clk_main_clk_clk                               : in  std_logic                     := 'X';             -- clk
			nios2_proc_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			sysid_qsys_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_proc_data_master_address                 : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_proc_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_proc_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_proc_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_proc_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_proc_data_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			nios2_proc_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_proc_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_proc_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_proc_instruction_master_address          : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_proc_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_proc_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_proc_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_proc_instruction_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			led_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                   : out std_logic;                                        -- write
			led_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                              : out std_logic;                                        -- chipselect
			nios2_proc_debug_mem_slave_address             : out std_logic_vector(8 downto 0);                     -- address
			nios2_proc_debug_mem_slave_write               : out std_logic;                                        -- write
			nios2_proc_debug_mem_slave_read                : out std_logic;                                        -- read
			nios2_proc_debug_mem_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_proc_debug_mem_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_proc_debug_mem_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_proc_debug_mem_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			nios2_proc_debug_mem_slave_debugaccess         : out std_logic;                                        -- debugaccess
			onchip_memory_s1_address                       : out std_logic_vector(21 downto 0);                    -- address
			onchip_memory_s1_write                         : out std_logic;                                        -- write
			onchip_memory_s1_read                          : out std_logic;                                        -- read
			onchip_memory_s1_readdata                      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			onchip_memory_s1_writedata                     : out std_logic_vector(63 downto 0);                    -- writedata
			onchip_memory_s1_byteenable                    : out std_logic_vector(7 downto 0);                     -- byteenable
			onchip_memory_s1_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			onchip_memory_s1_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			onchip_memory_s1_chipselect                    : out std_logic;                                        -- chipselect
			switcher_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			switcher_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_0_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component blinker_mm_interconnect_0;

	component blinker_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component blinker_irq_mapper;

	component blinker_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component blinker_rst_controller;

	component blinker_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component blinker_rst_controller_001;

	signal nios2_proc_debug_reset_request_reset                     : std_logic;                     -- nios2_proc:debug_reset_request -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_001:reset_in1]
	signal nios2_proc_data_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_proc_data_master_readdata -> nios2_proc:d_readdata
	signal nios2_proc_data_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:nios2_proc_data_master_waitrequest -> nios2_proc:d_waitrequest
	signal nios2_proc_data_master_debugaccess                       : std_logic;                     -- nios2_proc:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_proc_data_master_debugaccess
	signal nios2_proc_data_master_address                           : std_logic_vector(26 downto 0); -- nios2_proc:d_address -> mm_interconnect_0:nios2_proc_data_master_address
	signal nios2_proc_data_master_byteenable                        : std_logic_vector(3 downto 0);  -- nios2_proc:d_byteenable -> mm_interconnect_0:nios2_proc_data_master_byteenable
	signal nios2_proc_data_master_read                              : std_logic;                     -- nios2_proc:d_read -> mm_interconnect_0:nios2_proc_data_master_read
	signal nios2_proc_data_master_readdatavalid                     : std_logic;                     -- mm_interconnect_0:nios2_proc_data_master_readdatavalid -> nios2_proc:d_readdatavalid
	signal nios2_proc_data_master_write                             : std_logic;                     -- nios2_proc:d_write -> mm_interconnect_0:nios2_proc_data_master_write
	signal nios2_proc_data_master_writedata                         : std_logic_vector(31 downto 0); -- nios2_proc:d_writedata -> mm_interconnect_0:nios2_proc_data_master_writedata
	signal nios2_proc_instruction_master_readdata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_proc_instruction_master_readdata -> nios2_proc:i_readdata
	signal nios2_proc_instruction_master_waitrequest                : std_logic;                     -- mm_interconnect_0:nios2_proc_instruction_master_waitrequest -> nios2_proc:i_waitrequest
	signal nios2_proc_instruction_master_address                    : std_logic_vector(26 downto 0); -- nios2_proc:i_address -> mm_interconnect_0:nios2_proc_instruction_master_address
	signal nios2_proc_instruction_master_read                       : std_logic;                     -- nios2_proc:i_read -> mm_interconnect_0:nios2_proc_instruction_master_read
	signal nios2_proc_instruction_master_readdatavalid              : std_logic;                     -- mm_interconnect_0:nios2_proc_instruction_master_readdatavalid -> nios2_proc:i_readdatavalid
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata    : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_readdata    : std_logic_vector(31 downto 0); -- nios2_proc:debug_mem_slave_readdata -> mm_interconnect_0:nios2_proc_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_waitrequest : std_logic;                     -- nios2_proc:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_proc_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_debugaccess : std_logic;                     -- mm_interconnect_0:nios2_proc_debug_mem_slave_debugaccess -> nios2_proc:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_address     : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_proc_debug_mem_slave_address -> nios2_proc:debug_mem_slave_address
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_read        : std_logic;                     -- mm_interconnect_0:nios2_proc_debug_mem_slave_read -> nios2_proc:debug_mem_slave_read
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_proc_debug_mem_slave_byteenable -> nios2_proc:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_write       : std_logic;                     -- mm_interconnect_0:nios2_proc_debug_mem_slave_write -> nios2_proc:debug_mem_slave_write
	signal mm_interconnect_0_nios2_proc_debug_mem_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_proc_debug_mem_slave_writedata -> nios2_proc:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory_s1_chipselect            : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:az_cs
	signal mm_interconnect_0_onchip_memory_s1_readdata              : std_logic_vector(63 downto 0); -- onchip_memory:za_data -> mm_interconnect_0:onchip_memory_s1_readdata
	signal mm_interconnect_0_onchip_memory_s1_waitrequest           : std_logic;                     -- onchip_memory:za_waitrequest -> mm_interconnect_0:onchip_memory_s1_waitrequest
	signal mm_interconnect_0_onchip_memory_s1_address               : std_logic_vector(21 downto 0); -- mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:az_addr
	signal mm_interconnect_0_onchip_memory_s1_read                  : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_read -> mm_interconnect_0_onchip_memory_s1_read:in
	signal mm_interconnect_0_onchip_memory_s1_byteenable            : std_logic_vector(7 downto 0);  -- mm_interconnect_0:onchip_memory_s1_byteenable -> mm_interconnect_0_onchip_memory_s1_byteenable:in
	signal mm_interconnect_0_onchip_memory_s1_readdatavalid         : std_logic;                     -- onchip_memory:za_valid -> mm_interconnect_0:onchip_memory_s1_readdatavalid
	signal mm_interconnect_0_onchip_memory_s1_write                 : std_logic;                     -- mm_interconnect_0:onchip_memory_s1_write -> mm_interconnect_0_onchip_memory_s1_write:in
	signal mm_interconnect_0_onchip_memory_s1_writedata             : std_logic_vector(63 downto 0); -- mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:az_data
	signal mm_interconnect_0_switcher_s1_readdata                   : std_logic_vector(31 downto 0); -- switcher:readdata -> mm_interconnect_0:switcher_s1_readdata
	signal mm_interconnect_0_switcher_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switcher_s1_address -> switcher:address
	signal mm_interconnect_0_led_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_readdata                        : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_led_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_write                           : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal nios2_proc_irq_irq                                       : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_proc:irq
	signal rst_controller_reset_out_reset                           : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:sysid_qsys_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                       : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_proc_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                   : std_logic;                     -- rst_controller_001:reset_req -> [nios2_proc:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_onchip_memory_s1_read_ports_inv        : std_logic;                     -- mm_interconnect_0_onchip_memory_s1_read:inv -> onchip_memory:az_rd_n
	signal mm_interconnect_0_onchip_memory_s1_byteenable_ports_inv  : std_logic_vector(7 downto 0);  -- mm_interconnect_0_onchip_memory_s1_byteenable:inv -> onchip_memory:az_be_n
	signal mm_interconnect_0_onchip_memory_s1_write_ports_inv       : std_logic;                     -- mm_interconnect_0_onchip_memory_s1_write:inv -> onchip_memory:az_wr_n
	signal mm_interconnect_0_led_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal rst_controller_reset_out_reset_ports_inv                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [led:reset_n, onchip_memory:reset_n, switcher:reset_n, sysid_qsys_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv             : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> nios2_proc:reset_n

begin

	led : component blinker_led
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	nios2_proc : component blinker_nios2_proc
		port map (
			clk                                 => clk_clk,                                                  --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                   --                          .reset_req
			d_address                           => nios2_proc_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_proc_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_proc_data_master_read,                              --                          .read
			d_readdata                          => nios2_proc_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_proc_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_proc_data_master_write,                             --                          .write
			d_writedata                         => nios2_proc_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_proc_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_proc_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_proc_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_proc_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_proc_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_proc_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_proc_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_proc_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_proc_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_proc_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_proc_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_proc_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_proc_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_proc_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_proc_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_proc_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_proc_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	onchip_memory : component blinker_onchip_memory
		port map (
			clk            => clk_clk,                                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                -- reset.reset_n
			az_addr        => mm_interconnect_0_onchip_memory_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_onchip_memory_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_onchip_memory_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_onchip_memory_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_onchip_memory_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_onchip_memory_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_onchip_memory_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_onchip_memory_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_onchip_memory_s1_waitrequest,          --      .waitrequest
			zs_addr        => open,                                                    --  wire.export
			zs_ba          => open,                                                    --      .export
			zs_cas_n       => open,                                                    --      .export
			zs_cke         => open,                                                    --      .export
			zs_cs_n        => open,                                                    --      .export
			zs_dq          => open,                                                    --      .export
			zs_dqm         => open,                                                    --      .export
			zs_ras_n       => open,                                                    --      .export
			zs_we_n        => open                                                     --      .export
		);

	switcher : component blinker_switcher
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switcher_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_switcher_s1_readdata,   --                    .readdata
			in_port  => switcher_external_connection_export       -- external_connection.export
		);

	sysid_qsys_0 : component blinker_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component blinker_mm_interconnect_0
		port map (
			clk_main_clk_clk                               => clk_clk,                                                  --                             clk_main_clk.clk
			nios2_proc_reset_reset_bridge_in_reset_reset   => rst_controller_001_reset_out_reset,                       --   nios2_proc_reset_reset_bridge_in_reset.reset
			sysid_qsys_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                           -- sysid_qsys_0_reset_reset_bridge_in_reset.reset
			nios2_proc_data_master_address                 => nios2_proc_data_master_address,                           --                   nios2_proc_data_master.address
			nios2_proc_data_master_waitrequest             => nios2_proc_data_master_waitrequest,                       --                                         .waitrequest
			nios2_proc_data_master_byteenable              => nios2_proc_data_master_byteenable,                        --                                         .byteenable
			nios2_proc_data_master_read                    => nios2_proc_data_master_read,                              --                                         .read
			nios2_proc_data_master_readdata                => nios2_proc_data_master_readdata,                          --                                         .readdata
			nios2_proc_data_master_readdatavalid           => nios2_proc_data_master_readdatavalid,                     --                                         .readdatavalid
			nios2_proc_data_master_write                   => nios2_proc_data_master_write,                             --                                         .write
			nios2_proc_data_master_writedata               => nios2_proc_data_master_writedata,                         --                                         .writedata
			nios2_proc_data_master_debugaccess             => nios2_proc_data_master_debugaccess,                       --                                         .debugaccess
			nios2_proc_instruction_master_address          => nios2_proc_instruction_master_address,                    --            nios2_proc_instruction_master.address
			nios2_proc_instruction_master_waitrequest      => nios2_proc_instruction_master_waitrequest,                --                                         .waitrequest
			nios2_proc_instruction_master_read             => nios2_proc_instruction_master_read,                       --                                         .read
			nios2_proc_instruction_master_readdata         => nios2_proc_instruction_master_readdata,                   --                                         .readdata
			nios2_proc_instruction_master_readdatavalid    => nios2_proc_instruction_master_readdatavalid,              --                                         .readdatavalid
			led_s1_address                                 => mm_interconnect_0_led_s1_address,                         --                                   led_s1.address
			led_s1_write                                   => mm_interconnect_0_led_s1_write,                           --                                         .write
			led_s1_readdata                                => mm_interconnect_0_led_s1_readdata,                        --                                         .readdata
			led_s1_writedata                               => mm_interconnect_0_led_s1_writedata,                       --                                         .writedata
			led_s1_chipselect                              => mm_interconnect_0_led_s1_chipselect,                      --                                         .chipselect
			nios2_proc_debug_mem_slave_address             => mm_interconnect_0_nios2_proc_debug_mem_slave_address,     --               nios2_proc_debug_mem_slave.address
			nios2_proc_debug_mem_slave_write               => mm_interconnect_0_nios2_proc_debug_mem_slave_write,       --                                         .write
			nios2_proc_debug_mem_slave_read                => mm_interconnect_0_nios2_proc_debug_mem_slave_read,        --                                         .read
			nios2_proc_debug_mem_slave_readdata            => mm_interconnect_0_nios2_proc_debug_mem_slave_readdata,    --                                         .readdata
			nios2_proc_debug_mem_slave_writedata           => mm_interconnect_0_nios2_proc_debug_mem_slave_writedata,   --                                         .writedata
			nios2_proc_debug_mem_slave_byteenable          => mm_interconnect_0_nios2_proc_debug_mem_slave_byteenable,  --                                         .byteenable
			nios2_proc_debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_proc_debug_mem_slave_waitrequest, --                                         .waitrequest
			nios2_proc_debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_proc_debug_mem_slave_debugaccess, --                                         .debugaccess
			onchip_memory_s1_address                       => mm_interconnect_0_onchip_memory_s1_address,               --                         onchip_memory_s1.address
			onchip_memory_s1_write                         => mm_interconnect_0_onchip_memory_s1_write,                 --                                         .write
			onchip_memory_s1_read                          => mm_interconnect_0_onchip_memory_s1_read,                  --                                         .read
			onchip_memory_s1_readdata                      => mm_interconnect_0_onchip_memory_s1_readdata,              --                                         .readdata
			onchip_memory_s1_writedata                     => mm_interconnect_0_onchip_memory_s1_writedata,             --                                         .writedata
			onchip_memory_s1_byteenable                    => mm_interconnect_0_onchip_memory_s1_byteenable,            --                                         .byteenable
			onchip_memory_s1_readdatavalid                 => mm_interconnect_0_onchip_memory_s1_readdatavalid,         --                                         .readdatavalid
			onchip_memory_s1_waitrequest                   => mm_interconnect_0_onchip_memory_s1_waitrequest,           --                                         .waitrequest
			onchip_memory_s1_chipselect                    => mm_interconnect_0_onchip_memory_s1_chipselect,            --                                         .chipselect
			switcher_s1_address                            => mm_interconnect_0_switcher_s1_address,                    --                              switcher_s1.address
			switcher_s1_readdata                           => mm_interconnect_0_switcher_s1_readdata,                   --                                         .readdata
			sysid_qsys_0_control_slave_address             => mm_interconnect_0_sysid_qsys_0_control_slave_address,     --               sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata            => mm_interconnect_0_sysid_qsys_0_control_slave_readdata     --                                         .readdata
		);

	irq_mapper : component blinker_irq_mapper
		port map (
			clk        => clk_clk,                            --       clk.clk
			reset      => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sender_irq => nios2_proc_irq_irq                  --    sender.irq
		);

	rst_controller : component blinker_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_proc_debug_reset_request_reset, -- reset_in0.reset
			clk            => clk_clk,                              --       clk.clk
			reset_out      => rst_controller_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                 -- (terminated)
			reset_req_in0  => '0',                                  -- (terminated)
			reset_in1      => '0',                                  -- (terminated)
			reset_req_in1  => '0',                                  -- (terminated)
			reset_in2      => '0',                                  -- (terminated)
			reset_req_in2  => '0',                                  -- (terminated)
			reset_in3      => '0',                                  -- (terminated)
			reset_req_in3  => '0',                                  -- (terminated)
			reset_in4      => '0',                                  -- (terminated)
			reset_req_in4  => '0',                                  -- (terminated)
			reset_in5      => '0',                                  -- (terminated)
			reset_req_in5  => '0',                                  -- (terminated)
			reset_in6      => '0',                                  -- (terminated)
			reset_req_in6  => '0',                                  -- (terminated)
			reset_in7      => '0',                                  -- (terminated)
			reset_req_in7  => '0',                                  -- (terminated)
			reset_in8      => '0',                                  -- (terminated)
			reset_req_in8  => '0',                                  -- (terminated)
			reset_in9      => '0',                                  -- (terminated)
			reset_req_in9  => '0',                                  -- (terminated)
			reset_in10     => '0',                                  -- (terminated)
			reset_req_in10 => '0',                                  -- (terminated)
			reset_in11     => '0',                                  -- (terminated)
			reset_req_in11 => '0',                                  -- (terminated)
			reset_in12     => '0',                                  -- (terminated)
			reset_req_in12 => '0',                                  -- (terminated)
			reset_in13     => '0',                                  -- (terminated)
			reset_req_in13 => '0',                                  -- (terminated)
			reset_in14     => '0',                                  -- (terminated)
			reset_req_in14 => '0',                                  -- (terminated)
			reset_in15     => '0',                                  -- (terminated)
			reset_req_in15 => '0'                                   -- (terminated)
		);

	rst_controller_001 : component blinker_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_proc_debug_reset_request_reset,   -- reset_in0.reset
			reset_in1      => nios2_proc_debug_reset_request_reset,   -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	mm_interconnect_0_onchip_memory_s1_read_ports_inv <= not mm_interconnect_0_onchip_memory_s1_read;

	mm_interconnect_0_onchip_memory_s1_byteenable_ports_inv <= not mm_interconnect_0_onchip_memory_s1_byteenable;

	mm_interconnect_0_onchip_memory_s1_write_ports_inv <= not mm_interconnect_0_onchip_memory_s1_write;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of blinker
