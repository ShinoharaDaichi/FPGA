library verilog;
use verilog.vl_types.all;
entity add4bit_vlg_vec_tst is
end add4bit_vlg_vec_tst;
