library verilog;
use verilog.vl_types.all;
entity add1bit_vlg_vec_tst is
end add1bit_vlg_vec_tst;
