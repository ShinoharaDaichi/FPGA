library verilog;
use verilog.vl_types.all;
entity ex2 is
    port(
        x               : in     vl_logic;
        y               : in     vl_logic;
        f               : out    vl_logic
    );
end ex2;
