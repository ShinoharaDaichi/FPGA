library verilog;
use verilog.vl_types.all;
entity ex1I_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ex1I_vlg_check_tst;
