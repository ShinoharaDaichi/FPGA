library verilog;
use verilog.vl_types.all;
entity ex1I_vlg_vec_tst is
end ex1I_vlg_vec_tst;
