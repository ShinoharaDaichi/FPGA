library verilog;
use verilog.vl_types.all;
entity light2_vlg_vec_tst is
end light2_vlg_vec_tst;
