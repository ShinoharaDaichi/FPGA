
module test (
	clk_clk,
	reset_reset_n,
	spi_0_reset_reset_n);	

	input		clk_clk;
	input		reset_reset_n;
	input		spi_0_reset_reset_n;
endmodule
